`timescale 1ns / 1ps

module Sequence(
    input X,
    output reg Y,
    input CLK,
    input RST
);